library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;

entity InstructionMem is
	port(	PC :in std_logic_vector(15 downto 0);
			Instruction : out std_logic_vector(15 downto 0));
end InstructionMem;

architecture Fetch of InstructionMem is
	type ROM_arr_add is array (0 to 25) of std_logic_vector(15 downto 0);
	signal ROM : ROM_arr_add :=(
	"0100"&"001" & "000" &"000000",		--load Reg1
	"0100000000000000",		--load Reg0
	"0100010000000000",		--load Reg2
	"0100011000000000",		--load Reg3
	"0100100000000000",		--load Reg4
	"0100101000000000",		--load Reg5
	"0100110000000000",		--load Reg6
	
	"0110001011111110",		--load Reg1, Reg2, Reg3, Reg4, Reg5, Reg6
	
	"0001"&"001"&"010"&"000001",		--adi Reg2 = Reg1 + 1
	"0001010100011011",		--adi Reg4 = Reg2 + "011011"
	
	"0000010100011001",		--add Reg3 = Reg2 + Reg4
	
	"0011101000000011",		--lhi Reg5 = "11" & "0000000"
	
	"0101101010000001",		--store Reg5 into Memory location (Reg2 + 1) i.e., 2
	
	"0100110010000001",		--load Reg6 from Memory location (Reg2+1) i.e., 2
	
	"0111010011111111",		--SM
	
	"1000001000000010",		--jal PC to Reg1
	
	"1100100101111110",		--beq PC with "111110" if Reg4 = Reg5
	"1100101110000010", 		--beq PC with "000010" if Reg5 = Reg6
	
	"1111000000000000",		--unknown instruction
	
	"1001101100000000",		--jlr store PC to Reg5, branch PC to Reg4
	
	"0100001001000000",		--load Reg1
	"0100010001000000",		--load Reg2
	"0100011001000000",		--load Reg3
	"0100100001000000",		--load Reg4
	"0100101001000000",		--load Reg5
--	"0100110001000000",		--load Reg6
	
	
	
--	"0100001000000000",		--load Reg1 = 1
--	"0100010000000010",		--load Reg2 = 2
--	"0100011000000011",		--load Reg3 = 3
--	"0100100000000100",		--load Reg4 = 4
--	"0100101000000101",		--load Reg5 = 5
--	"0100110000000110",		--load Reg6 = 6
--	"0100111000000111",		--load Reg7 = 7
--	
--	"0000001010011001",		--add Reg3 = Reg1 + Reg2
--	"0000100101110010",		--add Reg6 = Reg4 + Reg5
--	
--	"0001001010000001",
--	"0001101110000001",
	
	
	
--"0100101000000001",
--"0100010000000010",
--"0100100000000011",
----"1000010000001000",
--"0010110110011000",
--"0000011011000001",
--
--"0000011011000001",
--"0001110000100010",
--"0000101101000001",
--"1001000000000011",

--								"0011"& "001"&"000000000",				--1
--								"0011"& "001"&"000000001",				--2
--								"0011"& "001"&"000000010",				--3
--								"0100"& "001"& "000"& "000001",
--								"0100"& "010"& "001"& "000001",
--								"0100"& "011"& "010"& "000001",
--								"0100"& "100"& "011"& "000001",
--								"0100"& "101"& "100"& "000001",
--								"0100"& "110"& "101"& "000001",
--								"0000"& "001"& "010"& "011"& "0"& "00",
--								
--								"0011"& "001"&"000000010",	
--								"0011"& "001"&"000000010",	
--								"0011"& "001"&"000000010",	
--								"0011"& "001"&"000000010",	
--								"0011"& "001"&"000000010",	
--								"0011"& "001"&"000000010",	
--								"0011"& "001"&"000000010",	
--								"0011"& "001"&"000000010",	
--								"0011"& "001"&"000000010",
--								"1001"& "001"&"000"&"000000",	
--								"0011"& "001"&"000000010"
"1111111000000000"	
								);

begin

	Instruction <= ROM(to_integer(unsigned(PC)));
		
end Fetch;

---------------------------------------------------------------------------------------------
